LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TOP IS
  
  PORT(
    A : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    B : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    CLK : IN STD_LOGIC;
    LOAD : IN STD_LOGIC;
    CLR : IN STD_LOGIC;
    END_F : OUT STD_LOGIC;
    Z : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)    
  );
  
END TOP;

ARCHITECTURE TOP_LEVEL OF TOP IS

-- PIPELINING THROUGH FLIP FLOP
COMPONENT DFF32 IS

  PORT(
     d : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
     sync_reset : IN STD_LOGIC;
     clk : IN STD_LOGIC;
     q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END COMPONENT;

COMPONENT DFF16 IS

  PORT(
     d : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
     sync_reset : IN STD_LOGIC;
     clk : IN STD_LOGIC;
     q : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END COMPONENT;

-- CONTROL & FLAGS THROUGH FLIP FLOP
COMPONENT DFF IS

    PORT(
	     d : IN STD_LOGIC;
       sync_reset : IN STD_LOGIC;
       clk : IN STD_LOGIC;
       q : OUT STD_LOGIC
     );
END COMPONENT;

-- EDGE TRIGGER 
COMPONENT EDGE_TRIG IS
  PORT(
    d : IN STD_LOGIC;
    clk : IN STD_LOGIC;
    edge : OUT STD_LOGIC
  );
END COMPONENT;

-- 16X16 MULTIPLIER
COMPONENT multi_16bit IS
  PORT (
    A : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    B : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    Z : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END COMPONENT;

SIGNAL A_IP, B_IP, A_REG, B_REG, STAGE1_B_Q : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL LD_POS, CLR_POS, LOAD_IN, FF0_LD_EN, FF0_CLR_EN : STD_LOGIC;
SIGNAL END_FLAG, CLR_FLAG, S0_EN_FF : STD_LOGIC;
SIGNAL PRODUCT_AB, S1_AxB : STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN
  A_IP <= ( 15 DOWNTO 0 => (NOT CLR)) AND A;
  B_IP <= ( 15 DOWNTO 0 => (NOT CLR)) AND B;
  
  FF0_POS_LD : EDGE_TRIG PORT MAP ( d => LOAD, clk => CLK, edge => LD_POS);
  FF0_POS_CLR : EDGE_TRIG PORT MAP ( d => CLR, clk => CLK, edge => CLR_POS);
    
 -- LOAD AT POS
 LOAD_IN <=  LD_POS OR CLR;
  
  -- LOAD INPUTS IN FLIP FLOP  
  FF0_A_IP : DFF16 PORT MAP ( d => A_IP, sync_reset => '0', clk => LOAD_IN, q => A_REG);
  FF0_B_IP : DFF16 PORT MAP ( d => B_IP, sync_reset => '0', clk => LOAD_IN, q => B_REG);
    
  -- END FLAG SETTING
  FF0_LD_EN <= CLK OR LD_POS;
  FF0_LD_EF: DFF PORT MAP  (d => LD_POS, sync_reset => '0', clk => FF0_LD_EN, q => END_FLAG);
    
  -- CLEAR FLAG SETTING
  FF0_CLR_EN <= CLR_POS;
  FF0_CLR_CF: DFF PORT MAP  (d => CLR, sync_reset => '0', clk => FF0_CLR_EN, q => CLR_FLAG);
    
  -- EQUATION STAGES 1/4[A x B]+1
  
  -- A x B USING 16BIT MULTIPLIER
  
  AB_MULTI_16 : multi_16bit PORT MAP (A => A_REG, B => B_REG, Z => PRODUCT_AB);
    
  S0_EN_FF <= END_FLAG OR CLR_FLAG;
  
  -- FLIP FLOP STAGE 1
  S1_AxB_FF : DFF32 PORT MAP (d => PRODUCT_AB, sync_reset => S0_EN_FF, clk => CLK, q => S1_AxB);
  
  

END TOP_LEVEL;