LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY DIV_BY_CONST IS
  GENERIC ( DIVISOR : INTEGER := 4);
  PORT(
    DIV : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    QUO : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
    
END DIV_BY_CONST;

ARCHITECTURE DIVISION OF DIV_BY_CONST IS
  
BEGIN
  
  --QUO <= CONV_STD_LOGIC_VECTOR((CONV_INTEGER(DIV)/DIVISOR),32);
  QUO <= "00" & DIV(31 DOWNTO 2);
  
END DIVISION;
