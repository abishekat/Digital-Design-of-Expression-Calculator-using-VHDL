LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY EDGE_TRIG IS
GENERIC (DELAY : TIME := 2 ns);
  PORT(
    d : IN STD_LOGIC;
    clk : IN STD_LOGIC;
    edge : OUT STD_LOGIC
  );
END EDGE_TRIG;
 
ARCHITECTURE EDGE_TRIGGER OF EDGE_TRIG IS
  
  SIGNAL regA, regB : STD_LOGIC;
  
BEGIN
	  regA <= d AFTER DELAY;
  EDT : PROCESS(d)
  
  BEGIN
	IF RISING_EDGE(clk) THEN
		edge <= d AND (NOT regA);
	END IF;
  END PROCESS;
  
END EDGE_TRIGGER;