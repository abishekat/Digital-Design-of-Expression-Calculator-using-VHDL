LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DFF IS

PORT(
	d : IN STD_LOGIC;
	enable : IN STD_LOGIC;
	clk : IN STD_LOGIC;
	q : OUT STD_LOGIC
);
END DFF;

ARCHITECTURE DFF_ARCH OF DFF IS
BEGIN

	PROCESS (clk, enable) IS
	BEGIN
	  IF FALLING_EDGE(clk) THEN
        IF (enable='1') THEN
          q <= d;
        ELSE
          q <= '0';
        END IF;
     END IF;
	END PROCESS;
END ARCHITECTURE DFF_ARCH;