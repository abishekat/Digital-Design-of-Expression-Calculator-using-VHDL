LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DIV_TB IS
END DIV_TB;

ARCHITECTURE TEST_BENCH OF DIV_TB IS

COMPONENT DIV_BY_CONST
PORT(
   DIV : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
   QUO : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
 );

END COMPONENT;

SIGNAL clk : STD_LOGIC := '0';
SIGNAL a, b : STD_LOGIC_VECTOR (31 DOWNTO 0);

CONSTANT clk_period : time := 10ns;

BEGIN
  uut: DIV_BY_CONST
  PORT MAP(
    DIV => a, QUO => b
  );
  
  
  PROCESS
  BEGIN
    clk <= '0';
    WAIT FOR clk_period/2;
    clk <= '1';
    WAIT FOR clk_period/2;
  
  END PROCESS;
  
  stimulus : PROCESS
  BEGIN
    a <= "00000000000000000000000000001000";
  WAIT FOR clk_period*2;
  a <= "00000000000000000000000000011000";
 WAIT FOR clk_period*3;
 a <= "00000000000000000000000000010000";
WAIT FOR  clk_period*4;
a <= "00000000000000000000000000001000";
WAIT FOR  clk_period*5;
a <= "00000000000000000000000000101000";
WAIT FOR  clk_period*6;
a <= "00000000000000000000000000100000";
WAIT FOR  clk_period*7;
a <= "00000000000000000000000010000000";
WAIT FOR  clk_period*8;
a <= "00000000000000000000000000000100";
WAIT FOR  clk_period*9;
a <= "00000000000000000000000100000000";
WAIT FOR  clk_period*10;
a <= "00000000000000000000000001000000";
WAIT FOR  clk_period*11;
  END PROCESS;

END TEST_BENCH;


