LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DFF32 IS


PORT(
  d : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
  sync_reset : IN STD_LOGIC;
  clk : IN STD_LOGIC;
  q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END DFF32;

ARCHITECTURE DFF_ARCH OF DFF32 IS
BEGIN

  PROCESS (clk, sync_reset) IS
  BEGIN
      IF(sync_reset='1') THEN
        q <= (OTHERS => '0');
      ELSIF(rising_edge(clk)) THEN
        q <= d;
      END IF;
  END PROCESS;
END ARCHITECTURE DFF_ARCH;