LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DIV_TB IS
END DIV_TB;

ARCHITECTURE TEST_BENCH OF DIV_TB IS

COMPONENT DIV_BY_CONST
PORT(
   DIV : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
   QUO : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
 );

END COMPONENT;

SIGNAL clk : STD_LOGIC := '0';
SIGNAL a, b : STD_LOGIC_VECTOR (31 DOWNTO 0);

CONSTANT clk_period : time := 10ns;

BEGIN
  uut: DIV_BY_CONST
  PORT MAP(
    DIV => a, QUO => b
  );
  
  
  PROCESS
  BEGIN
    clk <= '0';
    WAIT FOR clk_period/2;
    clk <= '1';
    WAIT FOR clk_period/2;
  
  END PROCESS;
  
  stimulus : PROCESS
  BEGIN
    a <= "00000000000000000000000000001000";
  WAIT;
  END PROCESS;

END TEST_BENCH;


