LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FA32_TB IS
END FA32_TB;

ARCHITECTURE TEST_BENCH OF FA32_TB IS

COMPONENT FullAdder32
PORT (
   A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
   B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
   Cin : IN STD_LOGIC;
   S : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
   Cout : OUT STD_LOGIC
 );

END COMPONENT;

SIGNAL clk, reset, cin, cout : STD_LOGIC := '0';
SIGNAL a, b, s : STD_LOGIC_VECTOR (31 DOWNTO 0);

CONSTANT clk_period : time := 10ns;

BEGIN
  uut: FullAdder32
  PORT MAP(
    A => a, B => b, Cin => cin, S => s, Cout => cout
  );
  
  
  PROCESS
  BEGIN
    clk <= '0';
    WAIT FOR clk_period/2;
    clk <= '1';
    WAIT FOR clk_period/2;
  
  END PROCESS;
  
  stimulus : PROCESS
  BEGIN
    a <= "00000000000000000000000000000001";
    b <= "00000000000000000000000000000010";
  WAIT;
  END PROCESS;

END TEST_BENCH;

