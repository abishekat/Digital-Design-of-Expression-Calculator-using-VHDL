LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TOP IS
  
  PORT(
    A : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    B : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    CLK : IN STD_LOGIC;
    LOAD : IN STD_LOGIC;
    CLR : IN STD_LOGIC;
    END_F : OUT STD_LOGIC;
    Z : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)    
  );
  
END TOP;

ARCHITECTURE TOP_LEVEL OF TOP IS

-- PIPELINING THROUGH FLIP FLOP
COMPONENT DFF32 IS

  PORT(
     d : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
     enable : IN STD_LOGIC;
     clk : IN STD_LOGIC;
     q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END COMPONENT;

COMPONENT DFF16 IS

  PORT(
     d : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
     enable : IN STD_LOGIC;
     clk : IN STD_LOGIC;
     q : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END COMPONENT;

-- CONTROL & FLAGS THROUGH FLIP FLOP
COMPONENT DFF IS

    PORT(
	     d : IN STD_LOGIC;
       enable : IN STD_LOGIC;
       clk : IN STD_LOGIC;
       q : OUT STD_LOGIC
     );
END COMPONENT;


-- 16X16 MULTIPLIER
COMPONENT multi_16bit IS
  PORT (
    X : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    Y : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    Z_P : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END COMPONENT;

COMPONENT FullAdder32
PORT (
   A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
   B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
   Cin : IN STD_LOGIC;
   S : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
   Cout : OUT STD_LOGIC
 );

END COMPONENT;

COMPONENT MUX2TO1 
  PORT(
    a : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    sel : IN STD_LOGIC;
    O: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END COMPONENT;

SIGNAL A_IP, B_IP, A_REG, B_REG : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL LD_POS, CLR_POS, LOAD_IN, FF0_LD_EN, FF0_CLR_EN, FA_32_COUT : STD_LOGIC;
SIGNAL END_FLAG, CLR_FLAG, S0_EN_FF, S1_END_FLAG, S1_CLR_FLAG, S1_EN_FF, S2_END_FLAG, S2_CLR_FLAG, S2_EN_FF  : STD_LOGIC;
SIGNAL PRODUCT_AB, S1_AxB: STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL S2_SR_DIV_VAL, S2_SR_OP, S3_ADD_OPERAND, Z_OUT, Z_REG  : STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN
  A_IP <= ( 15 DOWNTO 0 => (NOT CLR)) AND A;
  B_IP <= ( 15 DOWNTO 0 => (NOT CLR)) AND B;
    
 -- LOAD AT POS
 LD_POS <= LOAD;
 CLR_POS <= CLR;
 LOAD_IN <= LD_POS;
  
  -- LOAD INPUTS IN FLIP FLOP  
  FF0_A_IP : DFF16 PORT MAP ( d => A_IP, enable => LOAD_IN, clk => CLK, q => A_REG);
  FF0_B_IP : DFF16 PORT MAP ( d => B_IP, enable => LOAD_IN, clk => CLK, q => B_REG);
    
  -- END FLAG SETTING
  FF0_LD_EN <= CLK OR LD_POS;
  FF0_LD_EF: DFF PORT MAP  (d => LD_POS, enable => FF0_LD_EN, clk => CLK, q => END_FLAG);
    
  -- CLEAR FLAG SETTING
  FF0_CLR_EN <= CLR_POS;
  FF0_CLR_CF: DFF PORT MAP  (d => CLR, enable => FF0_CLR_EN, clk => CLK, q => CLR_FLAG);
    
  -- EQUATION STAGES 1/4[A x B]+1
  
  -- A x B USING 16BIT MULTIPLIER
  
  AB_MULTI_16 : multi_16bit PORT MAP (X => A_REG, Y => B_REG, Z_P => PRODUCT_AB);

  S0_EN_FF <= END_FLAG;
  
  -- FLIP FLOP STAGE 1
  S1_AxB_FF : DFF32 PORT MAP (d => PRODUCT_AB, enable => S0_EN_FF, clk => CLK, q => S1_AxB);
  S1_E_FLAG : DFF PORT MAP (d => END_FLAG, enable => END_FLAG, clk => CLK, q => S1_END_FLAG);
  S1_C_FLAG : DFF PORT MAP (d => CLR_FLAG, enable => CLR_FLAG, clk => CLK, q => S1_CLR_FLAG);
  
  S1_EN_FF <= S1_END_FLAG;
  
  --FLIP FLOP STAGE 2 (1/4 OPERATAION)
  S2_SR_DIV_VAL <= "00" & S1_AxB(31 DOWNTO 2);

  
  S2_SR_FF: DFF32 PORT MAP(d => S2_SR_DIV_VAL, enable => S1_EN_FF, clk => CLK, q => S2_SR_OP);
  S2_E_FLAG : DFF PORT MAP (d => S1_END_FLAG, enable => S1_END_FLAG, clk => CLK, q => S2_END_FLAG);
  S2_C_FLAG : DFF PORT MAP (d => S1_CLR_FLAG, enable => S1_CLR_FLAG, clk => CLK, q => S2_CLR_FLAG); 
  
  S2_EN_FF <= S2_END_FLAG;
  
  -- STAGE 3 ADDITION
  S3_ADD_OPERAND <= (0 => '1', OTHERS => '0');
  
  S3_ADD_FA : FullAdder32 PORT MAP (A => S2_SR_OP, B => S3_ADD_OPERAND, Cin => '0', S => Z_OUT, Cout => FA_32_COUT);
  
  MUX_OUT : MUX2TO1 PORT MAP (a => Z_OUT, b => (OTHERS => '0'), sel => S2_CLR_FLAG, O => Z_REG);
  
  Z <= Z_REG;  
  END_F <= S2_END_FLAG;
  
END TOP_LEVEL;
