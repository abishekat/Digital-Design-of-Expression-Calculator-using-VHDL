LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MUX2TO1 IS
  PORT(
    a : IN STD_LOGIC;
    b : IN STD_LOGIC;
    sel : IN STD_LOGIC;
    O: OUT STD_LOGIC
  );
END MUX2TO1;

ARCHITECTURE MUX OF MUX2TO1 IS

BEGIN
  PROCESS(a, b, sel)
    BEGIN
      IF sel = '0' then
        O <= a;
      ELSE
        O <= b;
      END IF;
    END PROCESS;

END MUX;