LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY EDGE_TRIG IS
  PORT(
    d : IN STD_LOGIC;
    clk : IN STD_LOGIC;
    edge : OUT STD_LOGIC
  );
END EDGE_TRIG;
 
ARCHITECTURE EDGE_TRIGGER OF EDGE_TRIG IS
  
  SIGNAL regA, regB : STD_LOGIC;
  
BEGIN
  EDT : PROCESS(clk)
  
  BEGIN
    IF rising_edge(clk) THEN
      regA <= d;
      regB <= regA;
    END IF;
  END PROCESS;
  
  edge <= regA AND (NOT regB);
  
END EDGE_TRIGGER;