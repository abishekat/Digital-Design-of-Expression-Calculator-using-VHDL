LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DFF IS

PORT(
	d : IN STD_LOGIC;
	sync_reset : IN STD_LOGIC;
	clk : IN STD_LOGIC;
	q : OUT STD_LOGIC
);
END DFF;

ARCHITECTURE DFF_ARCH OF DFF IS
BEGIN

	PROCESS (clk, sync_reset) IS
	BEGIN
			IF(sync_reset='1') THEN
				q <= '0';
			ELSIF(rising_edge(clk)) THEN
				q <= d;
			END IF;
	END PROCESS;
END ARCHITECTURE DFF_ARCH;