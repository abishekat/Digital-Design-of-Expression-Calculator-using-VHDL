LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY myAND IS
	PORT (
		a : IN STD_LOGIC;
		b : IN STD_LOGIC;
		Y : OUT STD_LOGIC
	);
END myAND;
ARCHITECTURE Behavioral OF myAND IS
BEGIN
	Y <= a AND b;
END Behavioral;